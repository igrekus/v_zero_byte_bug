module main

fn main() {
	// empty
}
