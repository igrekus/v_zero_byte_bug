module main
// empty
